library verilog;
use verilog.vl_types.all;
entity Adder_vlg_vec_tst is
end Adder_vlg_vec_tst;
