library verilog;
use verilog.vl_types.all;
entity CtrlLogic_vlg_vec_tst is
end CtrlLogic_vlg_vec_tst;
